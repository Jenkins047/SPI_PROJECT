send_data = 28'b0010110100111110001000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b1010110000010111101001000000;
expected_data = 28'b0000011100000000000000000000;

@(next_data);

send_data = 28'b1010001000000001001010000000;
expected_data = 28'b1111111111010000000000000000;

@(next_data);

send_data = 28'b0000011000100111100000000000;
expected_data = 28'b0000000000010000000000000000;

@(next_data);

send_data = 28'b0011111101011001100001000000;
expected_data = 28'b0101010100000000000000000000;

@(next_data);

send_data = 28'b0100011000001000000010000000;
expected_data = 28'b1000110001000000000000000000;

@(next_data);

send_data = 28'b0000110001011100100011000000;
expected_data = 28'b1010100101000000000000000000;

@(next_data);

send_data = 28'b0111111000110010000100000000;
expected_data = 28'b0000011000000000000000000000;

@(next_data);

send_data = 28'b0101001100001100100101000000;
expected_data = 28'b1111110001000000000000000000;

@(next_data);

send_data = 28'b1100110101111111000110000000;
expected_data = 28'b0111101000000000000000000000;

@(next_data);

send_data = 28'b0110100100111100000111000000;
expected_data = 28'b1011001101000000000000000000;

@(next_data);

send_data = 28'b1000011100010010101000000000;
expected_data = 28'b0000000000000000000000000000;

@(next_data);

send_data = 28'b0111000100111100001001000000;
expected_data = 28'b0000100100000000000000000000;

@(next_data);

send_data = 28'b1110100000110110001010000000;
expected_data = 28'b1111111111010000000000000000;

@(next_data);

send_data = 28'b1110011001100110000000000000;
expected_data = 28'b0000000000010000000000000000;

@(next_data);

send_data = 28'b0011011000111110100001000000;
expected_data = 28'b1011001001010000000000000000;

@(next_data);

send_data = 28'b1001110001101011100010000000;
expected_data = 28'b0100101100000000000000000000;

@(next_data);

send_data = 28'b0110011101110101100011000000;
expected_data = 28'b1011010001000000000000000000;

@(next_data);

send_data = 28'b1010101100110011000100000000;
expected_data = 28'b0011001100000000000000000000;

@(next_data);

send_data = 28'b0000011100011000100101000000;
expected_data = 28'b0101011000000000000000000000;

@(next_data);

send_data = 28'b0010101000011101000110000000;
expected_data = 28'b0000010000100000000000000000;

@(next_data);

send_data = 28'b1101011001000111100111000000;
expected_data = 28'b0010101000000000000000000000;

@(next_data);

send_data = 28'b0101010101001001001000000000;
expected_data = 28'b0000001000100000000000000000;

@(next_data);

send_data = 28'b0001110000010100101001000000;
expected_data = 28'b0000100100000000000000000000;

@(next_data);

send_data = 28'b0000101100100100001010000000;
expected_data = 28'b1111111111010000000000000000;

@(next_data);

send_data = 28'b0110010100010001000000000000;
expected_data = 28'b0000000000010000000000000000;

@(next_data);

send_data = 28'b1010101000011000100001000000;
expected_data = 28'b1000011101000000000000000000;

@(next_data);

send_data = 28'b1101001101100111100010000000;
expected_data = 28'b1001101101000000000000000000;

@(next_data);

send_data = 28'b1110011001001100000011000000;
expected_data = 28'b1110001101000000000000000000;

@(next_data);

send_data = 28'b0000000100010001000100000000;
expected_data = 28'b0111001100000000000000000000;

@(next_data);

send_data = 28'b1010000101110111000101000000;
expected_data = 28'b0000001000100000000000000000;

@(next_data);

send_data = 28'b1100001100111001000110000000;
expected_data = 28'b1111000101000000000000000000;

@(next_data);

send_data = 28'b1011110101100110000111000000;
expected_data = 28'b1011110101000000000000000000;

@(next_data);

send_data = 28'b0110010000110100001000000000;
expected_data = 28'b0000010000100000000000000000;

@(next_data);

send_data = 28'b1011111100111010101001000000;
expected_data = 28'b0000101000000000000000000000;

@(next_data);

send_data = 28'b1110101000111001001010000000;
expected_data = 28'b1111111111010000000000000000;

@(next_data);

send_data = 28'b1011110100111000000000000000;
expected_data = 28'b0000000000010000000000000000;

@(next_data);

send_data = 28'b1111011101110000000001000000;
expected_data = 28'b0010110100010000000000000000;

@(next_data);

send_data = 28'b1111101000001000000010000000;
expected_data = 28'b0001011100000000000000000000;

@(next_data);

send_data = 28'b1010111100101111100011000000;
expected_data = 28'b0001010100000000000000000000;

@(next_data);

send_data = 28'b0001000001001010100100000000;
expected_data = 28'b0101011100000000000000000000;

@(next_data);

send_data = 28'b0100010001110111000101000000;
expected_data = 28'b0010000000100000000000000000;

@(next_data);

send_data = 28'b0101101100111110000110000000;
expected_data = 28'b0110011000000000000000000000;

@(next_data);

send_data = 28'b0110110100011101100111000000;
expected_data = 28'b0101101100000000000000000000;

@(next_data);

send_data = 28'b0101101000100010101000000000;
expected_data = 28'b0000011100000000000000000000;

@(next_data);

send_data = 28'b0000010000100100001001000000;
expected_data = 28'b0000100100000000000000000000;

@(next_data);

send_data = 28'b1100000000011111101010000000;
expected_data = 28'b0000111100000000000000000000;

@(next_data);

send_data = 28'b0000000001101000100000000000;
expected_data = 28'b0000000000010000000000000000;

@(next_data);

send_data = 28'b0001001100101000000001000000;
expected_data = 28'b1101000101000000000000000000;

@(next_data);

send_data = 28'b0111001100010110100010000000;
expected_data = 28'b0100001100000000000000000000;

@(next_data);

send_data = 28'b0000010000001011000011000000;
expected_data = 28'b1010000101000000000000000000;

@(next_data);

send_data = 28'b0100000001011100100100000000;
expected_data = 28'b0000001000100000000000000000;

@(next_data);

send_data = 28'b1010101101000010100101000000;
expected_data = 28'b1000000001100000000000000000;

@(next_data);

send_data = 28'b0000111001010100000110000000;
expected_data = 28'b1111111001000000000000000000;

@(next_data);

send_data = 28'b0100110000010000100111000000;
expected_data = 28'b0000111000000000000000000000;

@(next_data);

send_data = 28'b1011010001011111101000000000;
expected_data = 28'b0000010000100000000000000000;

@(next_data);

send_data = 28'b0010101100100010101001000000;
expected_data = 28'b0000010100000000000000000000;

@(next_data);

send_data = 28'b0001110000111110101010000000;
expected_data = 28'b1111111111010000000000000000;

@(next_data);

expected_data = 28'b0000000000010000000000000000;