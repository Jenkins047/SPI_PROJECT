select_slave = 1;
send_request = 1;

send_data = 28'b1110001000011000100010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011000100110000011000000;
expected_data = 28'b0111000100000000000000000000;
@(next_data);

send_data = 28'b0001100101011000100100000000;
expected_data = 28'b1111101110100000000000000000;
@(next_data);

send_data = 28'b1110001100101010100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0011011100110010000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010001101101101000111000000;
expected_data = 28'b0110111010000000000000000000;
@(next_data);

send_data = 28'b1010010000111000001000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b0101000001111110101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001001001010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011101011101100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011111000101010000001000000;
expected_data = 28'b1100001010100000000000000000;
@(next_data);

send_data = 28'b1111001001100111100010000000;
expected_data = 28'b0111111000000000000000000000;
@(next_data);

send_data = 28'b1110011000100011000011000000;
expected_data = 28'b0111100110000000000000000000;
@(next_data);

send_data = 28'b0111010100101000000100000000;
expected_data = 28'b1011100110100000000000000000;
@(next_data);

send_data = 28'b0001010001001101100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0111101100001101100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101000011100100111000000;
expected_data = 28'b1111011000100000000000000000;
@(next_data);

send_data = 28'b1010100101001011001000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1010110001010100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000011000100101001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011010000111111000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100101000100111000001000000;
expected_data = 28'b1011001000100000000000000000;
@(next_data);

send_data = 28'b1100011100000010100010000000;
expected_data = 28'b0100111000000000000000000000;
@(next_data);

send_data = 28'b0001111000000000000011000000;
expected_data = 28'b0110001100000000000000000000;
@(next_data);

send_data = 28'b0010011100101000000100000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0011101000101110000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0001001101101101000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111010000100011100111000000;
expected_data = 28'b0010011010000000000000000000;
@(next_data);

send_data = 28'b1001000001011001001000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b1010001100100100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110001100111110001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001100001000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111101100010010000001000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b0011111000111110100010000000;
expected_data = 28'b0111111110000000000000000000;
@(next_data);

send_data = 28'b0010010100010100000011000000;
expected_data = 28'b0001111110000000000000000000;
@(next_data);

send_data = 28'b1001000000100001100100000000;
expected_data = 28'b1101111110100000000000000000;
@(next_data);

send_data = 28'b1100011000100011000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1001000100000011100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011111100001111000111000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b1101000001111001101000000000;
expected_data = 28'b0000010100000000000000000000;
@(next_data);

send_data = 28'b0010111001101101001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101000100001000101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001011100001100100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001010001010110100001000000;
expected_data = 28'b0011000000000000000000000000;
@(next_data);

send_data = 28'b1000110000101011000010000000;
expected_data = 28'b1011110100100000000000000000;
@(next_data);

send_data = 28'b1000110001010010000011000000;
expected_data = 28'b0100011010000000000000000000;
@(next_data);

send_data = 28'b1110100001010111100100000000;
expected_data = 28'b0111101100000000000000000000;
@(next_data);

send_data = 28'b1100011001011111000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1110001001000000000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110001000001010000111000000;
expected_data = 28'b1100010010100000000000000000;
@(next_data);

send_data = 28'b1011011000111111001000000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1101111000000111101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011001000110010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110100000011110100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111010100111101000001000000;
expected_data = 28'b1010010100100000000000000000;
@(next_data);

send_data = 28'b0011110100010101000010000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1111110001001001000011000000;
expected_data = 28'b0001111000000000000000000000;
@(next_data);

send_data = 28'b0011111000001010000100000000;
expected_data = 28'b0110111100000000000000000000;
@(next_data);

send_data = 28'b1101101101110000100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100011101001110100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010101101011011000111000000;
expected_data = 28'b1000111000100000000000000000;
@(next_data);

send_data = 28'b0110100000111000101000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b1101110000101010001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011110100100110101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101000001010100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001000101101000000001000000;
expected_data = 28'b1101111110100000000000000000;
@(next_data);

send_data = 28'b0011011100000101000010000000;
expected_data = 28'b1101000100100000000000000000;
@(next_data);

send_data = 28'b0011001100100101000011000000;
expected_data = 28'b0001101100000000000000000000;
@(next_data);

send_data = 28'b0111101001110101000100000000;
expected_data = 28'b1111110110100000000000000000;
@(next_data);

send_data = 28'b0100000101000011000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0101101100010111000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000000001100011000111000000;
expected_data = 28'b1011011010100000000000000000;
@(next_data);

send_data = 28'b1110001101110001001000000000;
expected_data = 28'b0000101110000000000000000000;
@(next_data);

send_data = 28'b1110101001100110001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000010000001011101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010010100011001100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111011101011000100001000000;
expected_data = 28'b1101100000100000000000000000;
@(next_data);

send_data = 28'b1011010100111111100010000000;
expected_data = 28'b1111011110100000000000000000;
@(next_data);

send_data = 28'b0000101100101101000011000000;
expected_data = 28'b0101101000000000000000000000;
@(next_data);

send_data = 28'b0101110001010001000100000000;
expected_data = 28'b1111010100100000000000000000;
@(next_data);

send_data = 28'b1100101100011100000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0001000100111100000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101111100100001100111000000;
expected_data = 28'b0010001000000000000000000000;
@(next_data);

send_data = 28'b1111111001110000001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0110000100101001101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110111101000011101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011101100010000100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101101101001000001000000;
expected_data = 28'b0101110000000000000000000000;
@(next_data);

send_data = 28'b0100110101000101000010000000;
expected_data = 28'b1101101100100000000000000000;
@(next_data);

send_data = 28'b0111001101000100000011000000;
expected_data = 28'b0010011010000000000000000000;
@(next_data);

send_data = 28'b0111101101010001100100000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1110010000011111100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1011001100011101000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101111100110000100111000000;
expected_data = 28'b0110011000000000000000000000;
@(next_data);

send_data = 28'b0110011000110111101000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b0011000100111101101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011111101101101001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010011000110000100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100101001010010100001000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b1110101101010001100010000000;
expected_data = 28'b1110111110100000000000000000;
@(next_data);

send_data = 28'b0111010101101001000011000000;
expected_data = 28'b0111010110000000000000000000;
@(next_data);

send_data = 28'b0100011100100110100100000000;
expected_data = 28'b1010111100100000000000000000;
@(next_data);

send_data = 28'b1001000001001011100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1110010101010110000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010110101000101100111000000;
expected_data = 28'b1100101000100000000000000000;
@(next_data);

send_data = 28'b1010000001000111001000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1110010001001000101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000110001100010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101011100110110100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100101000100111100001000000;
expected_data = 28'b0100010000000000000000000000;
@(next_data);

send_data = 28'b1101010001011101100010000000;
expected_data = 28'b0100111110000000000000000000;
@(next_data);

send_data = 28'b0010111100110111100011000000;
expected_data = 28'b0110101000000000000000000000;
@(next_data);

send_data = 28'b0000011101111100100100000000;
expected_data = 28'b1101000010100000000000000000;
@(next_data);

send_data = 28'b0110101001111011000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1010000000111110100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001000000110011100111000000;
expected_data = 28'b0100000010000000000000000000;
@(next_data);

send_data = 28'b0000101100011001101000000000;
expected_data = 28'b0000100100000000000000000000;
@(next_data);

send_data = 28'b1001110001001100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100100000111010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001100001011011000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011011101011000100001000000;
expected_data = 28'b0100111000000000000000000000;
@(next_data);

send_data = 28'b1010010000011110000010000000;
expected_data = 28'b1011011100100000000000000000;
@(next_data);

send_data = 28'b1101101101100111000011000000;
expected_data = 28'b0101001010000000000000000000;
@(next_data);

send_data = 28'b1101110001111010100100000000;
expected_data = 28'b0011010100000000000000000000;
@(next_data);

send_data = 28'b1010010101100100100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0011011101101001100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110011001101000000111000000;
expected_data = 28'b0110111010000000000000000000;
@(next_data);

send_data = 28'b1101101100100110001000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b0001000100100101101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011101001001000001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000110001010011100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001100000110001000001000000;
expected_data = 28'b0011001100000000000000000000;
@(next_data);

send_data = 28'b0101000100000011100010000000;
expected_data = 28'b0111101010000000000000000000;
@(next_data);

send_data = 28'b1100011101001010100011000000;
expected_data = 28'b0010100000000000000000000000;
@(next_data);

send_data = 28'b1011110101000101100100000000;
expected_data = 28'b0111101010000000000000000000;
@(next_data);

send_data = 28'b0000101100011010100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0101011000100111000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010010101101110000111000000;
expected_data = 28'b1010110000100000000000000000;
@(next_data);

send_data = 28'b0010000001011111001000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b1001010100001111001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000010000011000101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0010101101010001000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000100101011000100001000000;
expected_data = 28'b1100110110100000000000000000;
@(next_data);

send_data = 28'b0010011100111010000010000000;
expected_data = 28'b1011100110100000000000000000;
@(next_data);

send_data = 28'b0101111001010001000011000000;
expected_data = 28'b0001001110000000000000000000;
@(next_data);

send_data = 28'b0111101001111100100100000000;
expected_data = 28'b1111110110100000000000000000;
@(next_data);

send_data = 28'b0000000100001100000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1111111100000010000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101101101101011000111000000;
expected_data = 28'b1111111010100000000000000000;
@(next_data);

send_data = 28'b1011111000110100001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0001000000011110001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1001111101110111001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100011100000000100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011111101010011100001000000;
expected_data = 28'b1100100010100000000000000000;
@(next_data);

send_data = 28'b1100101000101010000010000000;
expected_data = 28'b1011111110100000000000000000;
@(next_data);

send_data = 28'b0001111000000101100011000000;
expected_data = 28'b0110010100000000000000000000;
@(next_data);

send_data = 28'b1011101000111100000100000000;
expected_data = 28'b1111010100100000000000000000;
@(next_data);

send_data = 28'b1000000100000100000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1000110001000010000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010111100100001100111000000;
expected_data = 28'b0001100000000000000000000000;
@(next_data);

send_data = 28'b0111001100010000001000000000;
expected_data = 28'b0000011110000000000000000000;
@(next_data);

send_data = 28'b0000010101000100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101101001101001101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000101000001010100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1000100000000000100001000000;
expected_data = 28'b1001111100100000000000000000;
@(next_data);

send_data = 28'b0011100001111000000010000000;
expected_data = 28'b1000100110100000000000000000;
@(next_data);

send_data = 28'b1010000000010000000011000000;
expected_data = 28'b0001110010000000000000000000;
@(next_data);

send_data = 28'b1111110100011100000100000000;
expected_data = 28'b1101111110100000000000000000;
@(next_data);

send_data = 28'b0001111100101001000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1011000101101010100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0101111001110000000111000000;
expected_data = 28'b0110001010000000000000000000;
@(next_data);

send_data = 28'b1101010001011001101000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1000110001001111101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110000000110011101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0111011000010100100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100100100011100000001000000;
expected_data = 28'b1001111100100000000000000000;
@(next_data);

send_data = 28'b1100010000000101000010000000;
expected_data = 28'b0111100110000000000000000000;
@(next_data);

send_data = 28'b1001010000110011000011000000;
expected_data = 28'b0110001010000000000000000000;
@(next_data);

send_data = 28'b1001101100110000100100000000;
expected_data = 28'b1111101110100000000000000000;
@(next_data);

send_data = 28'b0000011001111101100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0111100000111011100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100000001010000100111000000;
expected_data = 28'b1111000000100000000000000000;
@(next_data);

send_data = 28'b0101000101110100001000000000;
expected_data = 28'b0000110000000000000000000000;
@(next_data);

send_data = 28'b0101011001101001001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010111101010010101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110010000111111000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111111100111110000001000000;
expected_data = 28'b1110001000100000000000000000;
@(next_data);

send_data = 28'b0001110101101100100010000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1100001101001110000011000000;
expected_data = 28'b0000111010000000000000000000;
@(next_data);

send_data = 28'b1100001100001001000100000000;
expected_data = 28'b0111111110000000000000000000;
@(next_data);

send_data = 28'b1111100101100000100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0100001100101111100110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100001001011001000111000000;
expected_data = 28'b1000011010100000000000000000;
@(next_data);

send_data = 28'b0010110100111110001000000000;
expected_data = 28'b0000101000000000000000000000;
@(next_data);

send_data = 28'b1010110000010111101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010001000000001001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000011000100111100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011111101011001100001000000;
expected_data = 28'b0101010100000000000000000000;
@(next_data);

send_data = 28'b0100011000001000000010000000;
expected_data = 28'b1011111110100000000000000000;
@(next_data);

send_data = 28'b0000110001011100100011000000;
expected_data = 28'b0010001110000000000000000000;
@(next_data);

send_data = 28'b0111111000110010000100000000;
expected_data = 28'b1111011110100000000000000000;
@(next_data);

send_data = 28'b0101001100001100100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b1100110101111111000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110100100111100000111000000;
expected_data = 28'b1001101000100000000000000000;
@(next_data);

send_data = 28'b1000011100010010101000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b0111000100111100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110100000110110001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110011001100110000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0011011000111110100001000000;
expected_data = 28'b1011001000100000000000000000;
@(next_data);

send_data = 28'b1001110001101011100010000000;
expected_data = 28'b0111111110000000000000000000;
@(next_data);

send_data = 28'b0110011101110101100011000000;
expected_data = 28'b0100111000000000000000000000;
@(next_data);

send_data = 28'b1010101100110011000100000000;
expected_data = 28'b1001110000100000000000000000;
@(next_data);

send_data = 28'b0000011100011000100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0010101000011101000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101011001000111100111000000;
expected_data = 28'b0101010010000000000000000000;
@(next_data);

send_data = 28'b0101010101001001001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0001110000010100101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000101100100100001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110010100010001000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1010101000011000100001000000;
expected_data = 28'b1000011100100000000000000000;
@(next_data);

send_data = 28'b1101001101100111100010000000;
expected_data = 28'b1011101100100000000000000000;
@(next_data);

send_data = 28'b1110011001001100000011000000;
expected_data = 28'b0110100100000000000000000000;
@(next_data);

send_data = 28'b0000000100010001000100000000;
expected_data = 28'b0111111110000000000000000000;
@(next_data);

send_data = 28'b1010000101110111000101000000;
expected_data = 28'b0000001100000000000000000000;
@(next_data);

send_data = 28'b1100001100111001000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011110101100110000111000000;
expected_data = 28'b1000011010100000000000000000;
@(next_data);

send_data = 28'b0110010000110100001000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b1011111100111010101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1110101000111001001010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1011110100111000000000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1111011101110000000001000000;
expected_data = 28'b0010110100000000000000000000;
@(next_data);

send_data = 28'b1111101000001000000010000000;
expected_data = 28'b1111011110100000000000000000;
@(next_data);

send_data = 28'b1010111100101111100011000000;
expected_data = 28'b0111110100000000000000000000;
@(next_data);

send_data = 28'b0001000001001010100100000000;
expected_data = 28'b1111000000100000000000000000;
@(next_data);

send_data = 28'b0100010001110111000101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0101101100111110000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0110110100011101100111000000;
expected_data = 28'b1011011010100000000000000000;
@(next_data);

send_data = 28'b0101101000100010101000000000;
expected_data = 28'b0000011000000000000000000000;
@(next_data);

send_data = 28'b0000010000100100001001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100000000011111101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0000000001101000100000000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001001100101000000001000000;
expected_data = 28'b1101000100100000000000000000;
@(next_data);

send_data = 28'b0111001100010110100010000000;
expected_data = 28'b0101001100000000000000000000;
@(next_data);

send_data = 28'b0000010000001011000011000000;
expected_data = 28'b0011100100000000000000000000;
@(next_data);

send_data = 28'b0100000001011100100100000000;
expected_data = 28'b1111101110100000000000000000;
@(next_data);

send_data = 28'b1010101101000010100101000000;
expected_data = 28'b1111111100100000000000000000;
@(next_data);

send_data = 28'b0000111001010100000110000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100110000010000100111000000;
expected_data = 28'b0001110010000000000000000000;
@(next_data);

send_data = 28'b1011010001011111101000000000;
expected_data = 28'b0000101110000000000000000000;
@(next_data);

send_data = 28'b0010101100100010101001000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001110000111110101010000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);