select_slave = 0;
send_request = 1;

send_data = 20'b00011001101100010100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11100011010101010101;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b00110111011001000110;
expected_data = 20'b00000010000100000000;
@(next_data);

send_data = 20'b10100011110110100111;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b10100100011100001000;
expected_data = 20'b00001010001000000000;
@(next_data);

send_data = 20'b01010000111111011001;
expected_data = 20'b01010000001000000000;
@(next_data);

send_data = 20'b10110010100101011010;
expected_data = 20'b11001110100000000000;
@(next_data);

send_data = 20'b00000111101110110000;
expected_data = 20'b01001100000000000000;
@(next_data);

send_data = 20'b00111110010101000001;
expected_data = 20'b01101010001000000000;
@(next_data);

send_data = 20'b11110010110011110010;
expected_data = 20'b00111101000000000000;
@(next_data);

send_data = 20'b11100110010001100011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01110101010100000100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b00010100100110110101;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b01111011000110110110;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b11001010001110010111;
expected_data = 20'b00000001000100000000;
@(next_data);

send_data = 20'b10101001100101101000;
expected_data = 20'b00001000000100000000;
@(next_data);

send_data = 20'b10101100101010001001;
expected_data = 20'b11010100101000000000;
@(next_data);

send_data = 20'b10000110010010101010;
expected_data = 20'b11111010101000000000;
@(next_data);

send_data = 20'b00110100011111100000;
expected_data = 20'b10110110100000000000;
@(next_data);

send_data = 20'b01001010010011100001;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b11000111000001010010;
expected_data = 20'b11111010101000000000;
@(next_data);

send_data = 20'b00011110000000000011;
expected_data = 20'b00011110001000000000;
@(next_data);

send_data = 20'b00100111010100000100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b00111010010111000101;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b00010011110110100110;
expected_data = 20'b00000011001000000000;
@(next_data);

send_data = 20'b11110100010001110111;
expected_data = 20'b00000010000100000000;
@(next_data);

send_data = 20'b10010000101100101000;
expected_data = 20'b00001010001000000000;
@(next_data);

send_data = 20'b10100011010010001001;
expected_data = 20'b11011101101000000000;
@(next_data);

send_data = 20'b11100011011111001010;
expected_data = 20'b10011101100000000000;
@(next_data);

send_data = 20'b01000011000100000000;
expected_data = 20'b00110011001000000000;
@(next_data);

send_data = 20'b01111011001001000001;
expected_data = 20'b01011111001000000000;
@(next_data);

send_data = 20'b00111110011111010010;
expected_data = 20'b11000011101000000000;
@(next_data);

send_data = 20'b00100101001010000011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b10010000010000110100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11000110010001100101;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b10010001000001110110;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b10111111000111100111;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11010000111100111000;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b00101110110110101001;
expected_data = 20'b00101110001000000000;
@(next_data);

send_data = 20'b11010001000100011010;
expected_data = 20'b10101111101000000000;
@(next_data);

send_data = 20'b00010111000110010000;
expected_data = 20'b11111110100000000000;
@(next_data);

send_data = 20'b00010100101011010001;
expected_data = 20'b10111001100000000000;
@(next_data);

send_data = 20'b10001100010101100010;
expected_data = 20'b11111011100000000000;
@(next_data);

send_data = 20'b10001100101001000011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11101000101011110100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11000110101111100101;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b11100010100000000110;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11100010000101000111;
expected_data = 20'b00000001000100000000;
@(next_data);

send_data = 20'b10110110011111101000;
expected_data = 20'b00000101001000000000;
@(next_data);

send_data = 20'b11011110000011111001;
expected_data = 20'b10100010100000000000;
@(next_data);

send_data = 20'b10110010011001011010;
expected_data = 20'b11001110100000000000;
@(next_data);

send_data = 20'b01101000001111010000;
expected_data = 20'b00101011001000000000;
@(next_data);

send_data = 20'b11110101011110100001;
expected_data = 20'b10001111100000000000;
@(next_data);

send_data = 20'b00111101001010100010;
expected_data = 20'b11010111101000000000;
@(next_data);

send_data = 20'b11111100100100100011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b00111110000101000100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11011011111000010101;
expected_data = 20'b00000011001000000000;
@(next_data);

send_data = 20'b01000111100111010110;
expected_data = 20'b00000010000100000000;
@(next_data);

send_data = 20'b00101011101101100111;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01101000011100011000;
expected_data = 20'b00001001001000000000;
@(next_data);

send_data = 20'b11011100010101001001;
expected_data = 20'b10100100100000000000;
@(next_data);

send_data = 20'b00111101010011011010;
expected_data = 20'b00111101000000000000;
@(next_data);

send_data = 20'b11001010000101010000;
expected_data = 20'b10110101100000000000;
@(next_data);

send_data = 20'b10010001110100000001;
expected_data = 20'b01000001001000000000;
@(next_data);

send_data = 20'b00110111000010100010;
expected_data = 20'b11111101100000000000;
@(next_data);

send_data = 20'b00110011010010100011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01111010111010100100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01000001100001100101;
expected_data = 20'b00000110001000000000;
@(next_data);

send_data = 20'b01011011001011100110;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b10000000110001100111;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b11100011111000101000;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b11101010110011001001;
expected_data = 20'b10010110101000000000;
@(next_data);

send_data = 20'b10000100000101111010;
expected_data = 20'b11111100101000000000;
@(next_data);

send_data = 20'b10100101001100110000;
expected_data = 20'b01110010001000000000;
@(next_data);

send_data = 20'b11110111101100010001;
expected_data = 20'b01000110000000000000;
@(next_data);

send_data = 20'b10110101011111110010;
expected_data = 20'b11001010101000000000;
@(next_data);

send_data = 20'b00001011010110100011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01011100101000100100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11001011001110000101;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b00010001011110000110;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b11011111010000110111;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11111110111000001000;
expected_data = 20'b00000110001000000000;
@(next_data);

send_data = 20'b01100001010100111001;
expected_data = 20'b01100001000000000000;
@(next_data);

send_data = 20'b11101111100001111010;
expected_data = 20'b10010001100000000000;
@(next_data);

send_data = 20'b00111011001000010000;
expected_data = 20'b00011010000000000000;
@(next_data);

send_data = 20'b11001011110100100001;
expected_data = 20'b00011001000000000000;
@(next_data);

send_data = 20'b01001101100010100010;
expected_data = 20'b11110111100000000000;
@(next_data);

send_data = 20'b01110011100010000011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01111011101000110100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11100100001111110101;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b10110011001110100110;
expected_data = 20'b00000101001000000000;
@(next_data);

send_data = 20'b01011111011000010111;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01100110011011111000;
expected_data = 20'b00000110001000000000;
@(next_data);

send_data = 20'b00110001011110111001;
expected_data = 20'b00110001000000000000;
@(next_data);

send_data = 20'b00111111110110101010;
expected_data = 20'b00111111001000000000;
@(next_data);

send_data = 20'b10100110011000010000;
expected_data = 20'b01000101000000000000;
@(next_data);

send_data = 20'b01001010101001010001;
expected_data = 20'b11101111100000000000;
@(next_data);

send_data = 20'b11101011101000110010;
expected_data = 20'b01011100001000000000;
@(next_data);

send_data = 20'b01110101110100100011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01000111010011010100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b10010000100101110101;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b11100101101011000110;
expected_data = 20'b00000110001000000000;
@(next_data);

send_data = 20'b00101101100010110111;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b10100000100011101000;
expected_data = 20'b00001010001000000000;
@(next_data);

send_data = 20'b11100100100100011001;
expected_data = 20'b10011100101000000000;
@(next_data);

send_data = 20'b10001100110001011010;
expected_data = 20'b11110100100000000000;
@(next_data);

send_data = 20'b11010111011011010000;
expected_data = 20'b01101010001000000000;
@(next_data);

send_data = 20'b01001010010011110001;
expected_data = 20'b00000101001000000000;
@(next_data);

send_data = 20'b11010100101110110010;
expected_data = 20'b01101111001000000000;
@(next_data);

send_data = 20'b00101111011011110011;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b00000111111110010100;
expected_data = 20'b00000000001000000000;
@(next_data);

send_data = 20'b01101010111101100101;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b10100000011111010110;
expected_data = 20'b00000111000000000000;
@(next_data);

send_data = 20'b10010000011001110111;
expected_data = 20'b00000100000100000000;
@(next_data);

send_data = 20'b00001011001100111000;
expected_data = 20'b00001001001000000000;
@(next_data);

send_data = 20'b10011100100110001001;
expected_data = 20'b11100100101000000000;
@(next_data);

send_data = 20'b01001000011101011010;
expected_data = 20'b01001000001000000000;

@(next_data);
send_data = {8'd111, 8'd0, 4'd0};
expected_data = 20'b0000000000000000000000;
@(next_data);

send_data = {8'd99, 8'd203, 4'd0};
expected_data = {8'd111, 4'b0100, 9'b0};
@(next_data);

send_data = 20'b01100011110101010000;
expected_data = {8'b10001110, 4'b0100, 9'b0};
@(next_data);

send_data = 20'b10110011110000000000;
expected_data = 20'b0011100101000000000000;
@(next_data);

send_data = 20'b01110110011011110000;
expected_data = 20'b1100110101000000000000;
@(next_data);

send_data = 20'b10111100000100000001;
expected_data = 20'b0001110000000000000000;
@(next_data);

send_data = 20'b11011001001000010001;
expected_data = 20'b1011000101000000000000;
@(next_data);

send_data = 20'b10010011110100010001;
expected_data = 20'b1110000001000000000000;
@(next_data);

send_data = 20'b01001001000010010001;
expected_data = 20'b0000100100000000000000;
@(next_data);

send_data = 20'b10010001011111110010;
expected_data = 20'b0000001000000000000000;
@(next_data);

send_data = 20'b11111110111101110010;
expected_data = 20'b1011100101000000000000;
@(next_data);

send_data = 20'b01110101110111000010;
expected_data = 20'b0010010100000000000000;
@(next_data);

send_data = 20'b00010001001011000010;
expected_data = 20'b1010110001000000000000;
@(next_data);

send_data = 20'b10100010100111000011;
expected_data = 20'b1111110111000000000000;
@(next_data);

send_data = 20'b00111111000000010011;
expected_data = 20'b0000000100000000000000;
@(next_data);

send_data = 20'b01000100000000100011;
expected_data = 20'b1111100100000000000000;
@(next_data);

send_data = 20'b01001011000000110011;
expected_data = 20'b0100001000000000000000;
@(next_data);

send_data = 20'b01010101000000000100;
expected_data = 20'b0110000000000000000000;
@(next_data);

send_data = 20'b00001111000000010100;
expected_data = 20'b0101010100000000000000;
@(next_data);

send_data = 20'b11101011000000100100;
expected_data = 20'b0001110000000000000000;
@(next_data);

send_data = 20'b01001100000000110100;
expected_data = 20'b1110100100000000000000;
@(next_data);

send_data = 20'b00011001000000000101;
expected_data = 20'b0010010100000000000000;
@(next_data);

send_data = 20'b11000111011010110101;
expected_data = 20'b0000000100000000000000;
@(next_data);

send_data = 20'b11011011100001000101;
expected_data = 20'b0000011000000000000000;
@(next_data);

send_data = 20'b00101101101100110101;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00000001100111010111;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00010000111001100111;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00010000010111010111;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00100000000101010111;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00001000010000101000;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00110010001110001000;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00010110101011101000;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b01100111111100111000;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10000101011111111001;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b11010100010100101001;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b11110111101100111001;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10110100000010001001;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00101111011001101010;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10101101010001111010;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10011110000011011010;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b11010000110101101010;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b01001101010010001011;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10011001011010101011;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b01010100000100011011;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b11101011111100001011;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10011010101110101011;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10000010110010010101;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b10000010001010010110;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00010010011110110101;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00010010011010110110;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b11001011101001010101;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b11001011011101010110;
expected_data = 20'b0001001000000000000000;
@(next_data);

send_data = 20'b00110101111101100101;
expected_data = 20'b0001001000000000000000;
//@(next_data);

