select_slave = 0;
send_request = 1;

send_data = 28'b0110111100000000000000000000;
expected_data = 28'b0000000000000000000000000000;
@(next_data);

send_data = 28'b0110001101101010100000000000;
expected_data = 28'b0110111101000000000000000000;
@(next_data);

send_data = 28'b1011001101100000000000000000;
expected_data = 28'b1000111001010000000000000000;
@(next_data);

send_data = 28'b0111011000110111100000000000;
expected_data = 28'b1111001101010000000000000000;
@(next_data);

send_data = 28'b1011110000001000000001000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1101100100010000100001000000;
expected_data = 28'b1010110001010000000000000000;
@(next_data);

send_data = 28'b1001001101101000100001000000;
expected_data = 28'b1111100000010000000000000000;
@(next_data);

send_data = 28'b0100100100000100100001000000;
expected_data = 28'b0100001001000000000000000000;
@(next_data);

send_data = 28'b1001000100111111100010000000;
expected_data = 28'b0100000010000000000000000000;
@(next_data);

send_data = 28'b1111111001111011100010000000;
expected_data = 28'b1110111001010000000000000000;
@(next_data);

send_data = 28'b0111010101101110000010000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b0001000100010110000010000000;
expected_data = 28'b1010101100010000000000000000;
@(next_data);

send_data = 28'b1010001001001110000011000000;
expected_data = 28'b1111111101110000000000000000;
@(next_data);

send_data = 28'b0011111100000000100011000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0100010000000001000011000000;
expected_data = 28'b0111111001000000000000000000;
@(next_data);

send_data = 28'b0100101100000001100011000000;
expected_data = 28'b0001000010000000000000000000;
@(next_data);

send_data = 28'b0101010100000000000100000000;
expected_data = 28'b0101100000000000000000000000;
@(next_data);

send_data = 28'b0000111100000000100100000000;
expected_data = 28'b0101010101000000000000000000;
@(next_data);

send_data = 28'b1110101100000001000100000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0100110000000001100100000000;
expected_data = 28'b0011101001000000000000000000;
@(next_data);

send_data = 28'b0001100100000000000101000000;
expected_data = 28'b0000100101000000000000000000;
@(next_data);

send_data = 28'b1100011100110101100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1101101101000010000101000000;
expected_data = 28'b0000000110000000000000000000;
@(next_data);

send_data = 28'b0010110101011001100101000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b0000000101001110100111000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0001000001110011000111000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001000000101110100111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b0010000000001010100111000000;
expected_data = 28'b0000010010000000000000000000;
@(next_data);

send_data = 28'b0000100000100001001000000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b0011001000011100001000000000;
expected_data = 28'b0000110100000000000000000000;
@(next_data);

send_data = 28'b0001011001010111001000000000;
expected_data = 28'b0000101001000000000000000000;
@(next_data);

send_data = 28'b0110011101111001101000000000;
expected_data = 28'b0000100010000000000000000000;
@(next_data);

send_data = 28'b1000010100111111101001000000;
expected_data = 28'b0000010101000000000000000000;
@(next_data);

send_data = 28'b1101010000101001001001000000;
expected_data = 28'b1111101100010000000000000000;
@(next_data);

send_data = 28'b1111011101011001101001000000;
expected_data = 28'b1010110001010000000000000000;
@(next_data);

send_data = 28'b1011010000000100001001000000;
expected_data = 28'b1000100100010000000000000000;
@(next_data);

send_data = 28'b0010111100110011001010000000;
expected_data = 28'b1100110001010000000000000000;
@(next_data);

send_data = 28'b1010110100100011101010000000;
expected_data = 28'b0010111100000000000000000000;
@(next_data);

send_data = 28'b1001111000000110101010000000;
expected_data = 28'b1101001100010000000000000000;
@(next_data);

send_data = 28'b1101000001101011001010000000;
expected_data = 28'b1110001001010000000000000000;
@(next_data);

send_data = 28'b0100110100100100001011000000;
expected_data = 28'b1011000000010000000000000000;
@(next_data);

send_data = 28'b1001100100110101001011000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b0101010000001000101011000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1110101101111000001011000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1001101001011101001011000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1000001001100100100101000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b1000001000010100100110000000;
expected_data = 28'b0000001010000000000000000000;
@(next_data);

send_data = 28'b0001001000111101100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b0001001000110101100110000000;
expected_data = 28'b0000011001000000000000000000;
@(next_data);

send_data = 28'b1100101101010010100101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

send_data = 28'b1100101100111010100110000000;
expected_data = 28'b0000011100000000000000000000;
@(next_data);

send_data = 28'b0011010101111011000101000000;
expected_data = 28'b0000000001000000000000000000;
@(next_data);

