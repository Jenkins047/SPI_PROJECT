select_slave = 0;
send_request = 1;

send_data = {8'd111, 8'd0, 4'd0};
expected_data = 21'b0000000000000000000000;
@(next_data);

send_data = {8'd99, 8'd213, 4'd0};
expected_data = {8'd111, 4'b0100, 9'b0};
@(next_data);

send_data = 21'b01100011110101010000;
expected_data = {8'b10001110, 4'b0100, 9'b0};
@(next_data);

send_data = 21'b10110011110000000000;
expected_data = 21'b0011100101000000000000;
@(next_data);

send_data = 21'b01110110011011110000;
expected_data = 21'b1100110101000000000000;
@(next_data);

send_data = 21'b10111100000100000001;
expected_data = 21'b0001110000000000000000;
@(next_data);

send_data = 21'b11011001001000010001;
expected_data = 21'b1011000101000000000000;
@(next_data);

send_data = 21'b10010011110100010001;
expected_data = 21'b1110000001000000000000;
@(next_data);

send_data = 21'b01001001000010010001;
expected_data = 21'b0000100100000000000000;
@(next_data);

send_data = 21'b10010001011111110010;
expected_data = 21'b0000001000000000000000;
@(next_data);

send_data = 21'b11111110111101110010;
expected_data = 21'b1011100101000000000000;
@(next_data);

send_data = 21'b01110101110111000010;
expected_data = 21'b0010010100000000000000;
@(next_data);

send_data = 21'b00010001001011000010;
expected_data = 21'b1010110001000000000000;
@(next_data);

send_data = 21'b10100010100111000011;
expected_data = 21'b1111110111000000000000;
@(next_data);

send_data = 21'b00111111000000010011;
expected_data = 21'b0000000100000000000000;
@(next_data);

send_data = 21'b01000100000000100011;
expected_data = 21'b1111100100000000000000;
@(next_data);

send_data = 21'b01001011000000110011;
expected_data = 21'b0100001000000000000000;
@(next_data);

send_data = 21'b01010101000000000100;
expected_data = 21'b0110000000000000000000;
@(next_data);

send_data = 21'b00001111000000010100;
expected_data = 21'b0101010100000000000000;
@(next_data);

send_data = 21'b11101011000000100100;
expected_data = 21'b0001110000000000000000;
@(next_data);

send_data = 21'b01001100000000110100;
expected_data = 21'b1110100100000000000000;
@(next_data);

send_data = 21'b00011001000000000101;
expected_data = 21'b0010010100000000000000;
@(next_data);

send_data = 21'b11000111011010110101;
expected_data = 21'b0000000100000000000000;
@(next_data);

send_data = 21'b11011011100001000101;
expected_data = 21'b0000011000000000000000;
@(next_data);

send_data = 21'b00101101101100110101;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00000001100111010111;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00010000111001100111;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00010000010111010111;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00100000000101010111;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00001000010000101000;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00110010001110001000;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00010110101011101000;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b01100111111100111000;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10000101011111111001;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b11010100010100101001;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b11110111101100111001;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10110100000010001001;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00101111011001101010;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10101101010001111010;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10011110000011011010;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b11010000110101101010;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b01001101010010001011;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10011001011010101011;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b01010100000100011011;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b11101011111100001011;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10011010101110101011;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10000010110010010101;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b10000010001010010110;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00010010011110110101;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00010010011010110110;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b11001011101001010101;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b11001011011101010110;
expected_data = 21'b0001001000000000000000;
@(next_data);

send_data = 21'b00110101111101100101;
expected_data = 21'b0001001000000000000000;
@(next_data);